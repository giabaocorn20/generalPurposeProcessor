library verilog;
use verilog.vl_types.all;
entity lab6_vlg_vec_tst is
end lab6_vlg_vec_tst;
